<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-98.4076,24.3287,186.779,-116.634</PageViewport>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>39.5,-5.5</position>
<gparam>LABEL_TEXT NOR Gate As UNIVERSAL</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>56.5,-23</position>
<gparam>LABEL_TEXT AND GATE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>39.5,-29</position>
<gparam>LABEL_TEXT -------------------------------------------------------------------------</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>BE_NOR2</type>
<position>38,-35</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>28,-33</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>28,-37</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>BE_NOR2</type>
<position>47,-35</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>GA_LED</type>
<position>53,-35</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>58.5,-35</position>
<gparam>LABEL_TEXT OR GATE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>39.5,-40</position>
<gparam>LABEL_TEXT -------------------------------------------------------------------------</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>41.5,-83</position>
<gparam>LABEL_TEXT --------------------------------------------------------------------</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>BE_NOR2</type>
<position>37,-12</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_TOGGLE</type>
<position>29,-12</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>83</ID>
<type>GA_LED</type>
<position>44,-12</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>50.5,-12</position>
<gparam>LABEL_TEXT NOT GATE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>26.5,-11.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>39.5,-15.5</position>
<gparam>LABEL_TEXT -------------------------------------------------------------------------</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>BE_NOR2</type>
<position>37,-20</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>90</ID>
<type>BE_NOR2</type>
<position>37,-26</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_TOGGLE</type>
<position>28,-20</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_TOGGLE</type>
<position>28,-26</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>93</ID>
<type>BE_NOR2</type>
<position>45,-23</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>GA_LED</type>
<position>51,-23</position>
<input>
<ID>N_in0</ID>49 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>25.5,-19.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>25.5,-26</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-34,32.5,-33</points>
<intersection>-34 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-33,32.5,-33</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-34,35,-34</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-37,32.5,-36</points>
<intersection>-37 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-37,32.5,-37</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-36,35,-36</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-36,42.5,-34</points>
<intersection>-36 3</intersection>
<intersection>-35 1</intersection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-35,42.5,-35</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-34,44,-34</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>42.5,-36,44,-36</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-35,52,-35</points>
<connection>
<GID>9</GID>
<name>N_in0</name></connection>
<connection>
<GID>7</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-13,32.5,-11</points>
<intersection>-13 3</intersection>
<intersection>-12 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-12,32.5,-12</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-11,34,-11</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32.5,-13,34,-13</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-12,43,-12</points>
<connection>
<GID>83</GID>
<name>N_in0</name></connection>
<connection>
<GID>79</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-21,32.5,-19</points>
<intersection>-21 3</intersection>
<intersection>-20 4</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-19,34,-19</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32.5,-21,34,-21</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>30,-20,32.5,-20</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-27,32.5,-25</points>
<intersection>-27 3</intersection>
<intersection>-26 4</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-25,34,-25</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32.5,-27,34,-27</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>30,-26,32.5,-26</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-22,41,-20</points>
<intersection>-22 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-22,42,-22</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-20,41,-20</points>
<connection>
<GID>89</GID>
<name>OUT</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-26,41,-24</points>
<intersection>-26 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-24,42,-24</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-26,41,-26</points>
<connection>
<GID>90</GID>
<name>OUT</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-23,50,-23</points>
<connection>
<GID>94</GID>
<name>N_in0</name></connection>
<connection>
<GID>93</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 1>
<page 2>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 2>
<page 3>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 3>
<page 4>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 4>
<page 5>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 5>
<page 6>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 6>
<page 7>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 7>
<page 8>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 8>
<page 9>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 9></circuit>