<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-48,51,74.4,-9.5</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>-20,44</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>-29.5,46</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>-29.5,42</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>-13.5,44</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AE_OR2</type>
<position>-20,35</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>-29.5,36.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>-29.5,33</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>-13,35</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AE_SMALL_INVERTER</type>
<position>-20,28</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>-29.5,28</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>-13,28</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AI_XOR2</type>
<position>-19.5,21</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>-13,21</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>-29.5,22.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>-29.5,19.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>0,44.5</position>
<gparam>LABEL_TEXT AND GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>-1.5,35.5</position>
<gparam>LABEL_TEXT OR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>-0.5,28.5</position>
<gparam>LABEL_TEXT NOT GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AO_XNOR2</type>
<position>-19.5,12.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>GA_LED</type>
<position>-13,12.5</position>
<input>
<ID>N_in0</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>-30,14</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>-30,11</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>0.5,21.5</position>
<gparam>LABEL_TEXT EXOR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>1.5,13</position>
<gparam>LABEL_TEXT EXNOR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>BE_NOR2</type>
<position>-19.5,5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>-30,6.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>-30,3.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>GA_LED</type>
<position>-13,5</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>-0.5,5.5</position>
<gparam>LABEL_TEXT NOR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>BA_NAND2</type>
<position>-19,-2.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>-30,-1</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>-30,-4</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>60</ID>
<type>GA_LED</type>
<position>-12,-2.5</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>1,-2</position>
<gparam>LABEL_TEXT NAND GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27.5,46,-23,46</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-23 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-23,45,-23,46</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>46 1</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27.5,42,-23,42</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-23 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-23,42,-23,43</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>42 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17,44,-14.5,44</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>14</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,36,-25,36.5</points>
<intersection>36 1</intersection>
<intersection>36.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,36,-23,36</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27.5,36.5,-25,36.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,33,-25,34</points>
<intersection>33 2</intersection>
<intersection>34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,34,-23,34</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27.5,33,-25,33</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17,35,-14,35</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<connection>
<GID>16</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27.5,28,-22,28</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-18,28,-14,28</points>
<connection>
<GID>28</GID>
<name>N_in0</name></connection>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16.5,21,-14,21</points>
<connection>
<GID>32</GID>
<name>N_in0</name></connection>
<connection>
<GID>30</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,22,-25,22.5</points>
<intersection>22 1</intersection>
<intersection>22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,22,-22.5,22</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27.5,22.5,-25,22.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,19.5,-25,20</points>
<intersection>19.5 2</intersection>
<intersection>20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,20,-22.5,20</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27.5,19.5,-25,19.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,13.5,-25,14</points>
<intersection>13.5 1</intersection>
<intersection>14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,13.5,-22.5,13.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28,14,-25,14</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,11,-25,11.5</points>
<intersection>11 2</intersection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,11.5,-22.5,11.5</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28,11,-25,11</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16.5,12.5,-14,12.5</points>
<connection>
<GID>43</GID>
<name>N_in0</name></connection>
<connection>
<GID>42</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16.5,5,-14,5</points>
<connection>
<GID>52</GID>
<name>N_in0</name></connection>
<connection>
<GID>49</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,6,-25,6.5</points>
<intersection>6 1</intersection>
<intersection>6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,6,-22.5,6</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28,6.5,-25,6.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,3.5,-25,4</points>
<intersection>3.5 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,4,-22.5,4</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28,3.5,-25,3.5</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16,-2.5,-13,-2.5</points>
<connection>
<GID>60</GID>
<name>N_in0</name></connection>
<connection>
<GID>55</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,-4,-25,-3.5</points>
<intersection>-4 2</intersection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,-3.5,-22,-3.5</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28,-4,-25,-4</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,-1.5,-25,-1</points>
<intersection>-1.5 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,-1.5,-22,-1.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28,-1,-25,-1</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>